library verilog;
use verilog.vl_types.all;
entity vrf_timer_1s is
end vrf_timer_1s;
