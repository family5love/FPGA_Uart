library verilog;
use verilog.vl_types.all;
entity uart_rxd_vrf is
end uart_rxd_vrf;
